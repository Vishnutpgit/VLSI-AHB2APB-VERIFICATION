package bus_pkg ;
 
  import uvm_pkg::*;

`include "uvm_macros.svh" 
`include "mst_agt_config.sv"
`include "slv_agt_config.sv"
`include "env_config.sv"

`include "write_xtn.sv"
`include "read_xtn.sv"
`include "slv_monitor.sv"
`include "slv_driver.sv"
`include "slv_sequencer.sv"
`include "slv_agt.sv"
`include "slv_sequence.sv"

`include "mst_monitor.sv"
`include "mst_driver.sv"
`include "mst_sequencer.sv"
`include "mst_agt.sv"
`include "mst_sequence.sv"

`include "sb.sv"

`include "env.sv"
`include "test.sv"

endpackage
